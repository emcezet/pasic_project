`define SYMBOL_W 8
`define SYMBOL_NUM 8
`define DATA_W 8
`define TID_W 8
`define TDEST_W 8
`define TUSER_W 8

`define NUM_PORTS 4
`define PORT_WIDTH 128
`define FIFO_DEPTH 16
`define LOCAL_ADR 0

